library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity led_blinker_tb is
end led_blinker_tb;
component led_blinker_tb is
    port (

	 )
