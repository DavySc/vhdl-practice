library ieee;
use ieee.std_logic_1164.all;

entity alu4 is
	port(
	        
	    )
